----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:59:29 04/13/2016 
-- Design Name: 
-- Module Name:    delete - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity delete is
	port (
		inp : in std_logic_vector(4 downto 0):=(others=>'0');
		outp : out std_logic_vector(2 downto 0):=(others=>'0')
	);
end delete;

architecture Behavioral of delete is

begin
		outp <= inp(2 downto 0);


end Behavioral;

